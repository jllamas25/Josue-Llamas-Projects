`timescale 1ns / 1ps

module Or16bit(s,a,b);
    input [15:0] a,b;
    output [15:0] s;
    
	 or g[15:0] ( s,a,b);





endmodule
